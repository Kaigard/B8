module testRom (
    input logic clk,
    input logic reset_n,
    input logic request_i,
    input logic [31:0] instAddr_i,
    output logic [31:0] inst_o,
    output logic dataOk_o
);

    reg [7:0] romReg [10'h3FF * 4 : 0];

    initial begin
        $readmemh("code.mem", romReg);
    end

    /*
    always @(posedge clk or negedge reset_n) begin
        if(~reset_n) begin
            inst_o <= 32'b0;
            dataOk_o <= 1'b0;
        end else if(request_i) begin
            inst_o <= {romReg[instAddr_i], romReg[instAddr_i + 1], romReg[instAddr_i + 2], romReg[instAddr_i + 3]};
            dataOk_o <= 1'b1;
        end else begin
            dataOk_o <= 1'b0;
        end
    end
    */
    
    assign dataOk_o = 1'b1;
    assign inst_o = {romReg[instAddr_i], romReg[instAddr_i + 1], romReg[instAddr_i + 2], romReg[instAddr_i + 3]};
     
endmodule