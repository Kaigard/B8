`define TestMode 1
module BnineCore (
    input clk,
    input reset_n,
    //For Test
    input jumpFlag_i,
    input [31:0] jumpAddr_i,
    input ready_test
);

    wire way0_dataOk_i;
    wire way0_request_o;
    wire way1_dataOk_i;
    wire way1_request_o;
    wire [31:0] way0_inst_fetch_i;
    wire [31:0] way0_instAddr_fetch_o;
    wire [31:0] way1_inst_fetch_i;
    wire [31:0] way1_instAddr_fetch_o;

    testRom u_testRom_way0 (
        .clk(clk),
        .reset_n(reset_n),
        .request_i(way0_request_o),
        .instAddr_i(way0_instAddr_fetch_o),
        .inst_o(way0_inst_fetch_i),
        .dataOk_o(way0_dataOk_i)
    );

    testRom u_testRom_way1 (
        .clk(clk),
        .reset_n(reset_n),
        .request_i(way1_request_o),
        .instAddr_i(way1_instAddr_fetch_o),
        .inst_o(way1_inst_fetch_i),
        .dataOk_o(way1_dataOk_i)
    );

    BnineCore_way0 B_BnineCore_way0(
        .clk(clk),
        .reset_n(reset_n),
        .way0_dataOk_i(way0_dataOk_i),
        .way0_inst_fetch_i(way0_inst_fetch_i),
        .way0_request_o(way0_request_o),
        .way0_instAddr_fetch_o(way0_instAddr_fetch_o),
        // For Test
        .jumpFlag_i(jumpFlag_i),
        .jumpAddr_i(jumpAddr_i),
        .ready_test(ready_test)
    );

    BnineCore_way1 B_BnineCore_way1(
        .clk(clk),
        .reset_n(reset_n),
        .way1_dataOk_i(way1_dataOk_i),
        .way1_inst_fetch_i(way1_inst_fetch_i),
        .way1_request_o(way1_request_o),
        .way1_instAddr_fetch_o(way1_instAddr_fetch_o),
        // For Test
        .jumpFlag_i(jumpFlag_i),
        .jumpAddr_i(jumpAddr_i),
        .ready_test(ready_test)
    );

endmodule