module ExecuteUnit_way0(
    

);


endmodule